`define DELAY 20
module nine_to_one_mux_testbench ();

reg [5:0] funct;
reg [31:0] sll_out, srl_out, sra_out, add_out, addu_out, and_out, or_out, sub_out, sltu_out;
wire [31:0] out;

nine_to_one_mux muxtb(funct, sll_out, srl_out, sra_out, add_out, addu_out, and_out, or_out, sub_out, sltu_out, out);

initial begin
	  /*
	  6'b000000 : out = sll_out;
	  6'b000010 : out = srl_out;
	  6'b000011 : out = sra_out;
	  6'b100000 : out = add_out;
	  6'b100001 : out = addu_out;
	  6'b100100 : out = and_out;
	  6'b100101 : out = or_out;
	  6'b100010 : out = sub_out;
	  6'b101011 : out = sltu_out;
	*/
sll_out  = 32'b00000000000000000000000000000000;
srl_out  = 32'b00000000000000000000000000000001;
sra_out  = 32'b00000000000000000000000000000010;
add_out  = 32'b00000000000000000000000000000011;
addu_out = 32'b00000000000000000000000000000100;
and_out  = 32'b00000000000000000000000000000101;
or_out   = 32'b00000000000000000000000000000110;
sub_out  = 32'b00000000000000000000000000000111;
sltu_out = 32'b00000000000000000000000000001000;
funct    =  6'b000000;
#`DELAY;
sll_out  = 32'b00000000000000000000000000000000;
srl_out  = 32'b00000000000000000000000000000001;
sra_out  = 32'b00000000000000000000000000000010;
add_out  = 32'b00000000000000000000000000000011;
addu_out = 32'b00000000000000000000000000000100;
and_out  = 32'b00000000000000000000000000000101;
or_out   = 32'b00000000000000000000000000000110;
sub_out  = 32'b00000000000000000000000000000111;
sltu_out = 32'b00000000000000000000000000001000;
funct    =  6'b100001;
#`DELAY;
sll_out  = 32'b00000000000000000000000000000000;
srl_out  = 32'b00000000000000000000000000000001;
sra_out  = 32'b00000000000000000000000000000010;
add_out  = 32'b00000000000000000000000000000011;
addu_out = 32'b00000000000000000000000000000100;
and_out  = 32'b00000000000000000000000000000101;
or_out   = 32'b00000000000000000000000000000110;
sub_out  = 32'b00000000000000000000000000000111;
sltu_out = 32'b00000000000000000000000000001000;
funct    =  6'b100100;
#`DELAY;

end


initial
begin
$monitor("%6b     \n%32b \n\n", funct, out);
end
 
endmodule
